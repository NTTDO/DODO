module DEQAM(
	input [63:0] data_in,
	output reg [5:0] data_out
);
	always @(*) begin
		case(data_in)
64'b1100000011100000000000000000000001000000111000000000000000000000: data_out = 6'b000000;
64'b1100000010100000000000000000000001000000111000000000000000000000: data_out = 6'b000001;
64'b1100000001000000000000000000000001000000111000000000000000000000: data_out = 6'b000011;
64'b1011111110000000000000000000000001000000111000000000000000000000: data_out = 6'b000010;
64'b0011111110000000000000000000000001000000111000000000000000000000: data_out = 6'b000110;
64'b0100000001000000000000000000000001000000111000000000000000000000: data_out = 6'b000111;
64'b0100000010100000000000000000000001000000111000000000000000000000: data_out = 6'b000101;
64'b0100000011100000000000000000000001000000111000000000000000000000: data_out = 6'b000100;
64'b0100000011100000000000000000000001000000101000000000000000000000: data_out = 6'b001100;
64'b0100000010100000000000000000000001000000101000000000000000000000: data_out = 6'b001101;
64'b0100000001000000000000000000000001000000101000000000000000000000: data_out = 6'b001111;
64'b0011111110000000000000000000000001000000101000000000000000000000: data_out = 6'b001110;
64'b1011111110000000000000000000000001000000101000000000000000000000: data_out = 6'b001010;
64'b1100000001000000000000000000000001000000101000000000000000000000: data_out = 6'b001011;
64'b1100000010100000000000000000000001000000101000000000000000000000: data_out = 6'b001001;
64'b1100000011100000000000000000000001000000101000000000000000000000: data_out = 6'b001000;
64'b1100000011100000000000000000000001000000010000000000000000000000: data_out = 6'b011000;
64'b1100000010100000000000000000000001000000010000000000000000000000: data_out = 6'b011001;
64'b1100000001000000000000000000000001000000010000000000000000000000: data_out = 6'b011011;
64'b1011111110000000000000000000000001000000010000000000000000000000: data_out = 6'b011010;
64'b0011111110000000000000000000000001000000010000000000000000000000: data_out = 6'b011110;
64'b0100000001000000000000000000000001000000010000000000000000000000: data_out = 6'b011111;
64'b0100000010100000000000000000000001000000010000000000000000000000: data_out = 6'b011101;
64'b0100000011100000000000000000000001000000010000000000000000000000: data_out = 6'b011100;
64'b0100000011100000000000000000000000111111100000000000000000000000: data_out = 6'b010100;
64'b0100000010100000000000000000000000111111100000000000000000000000: data_out = 6'b010101;
64'b0100000001000000000000000000000000111111100000000000000000000000: data_out = 6'b010111;
64'b0011111110000000000000000000000000111111100000000000000000000000: data_out = 6'b010110;
64'b1011111110000000000000000000000000111111100000000000000000000000: data_out = 6'b010010;
64'b1100000001000000000000000000000000111111100000000000000000000000: data_out = 6'b010011;
64'b1100000010100000000000000000000000111111100000000000000000000000: data_out = 6'b010001;
64'b1100000011100000000000000000000000111111100000000000000000000000: data_out = 6'b010000;
64'b1100000011100000000000000000000010111111100000000000000000000000: data_out = 6'b110000;
64'b1100000010100000000000000000000010111111100000000000000000000000: data_out = 6'b110001;
64'b1100000001000000000000000000000010111111100000000000000000000000: data_out = 6'b110011;
64'b1011111110000000000000000000000010111111100000000000000000000000: data_out = 6'b110010;
64'b0011111110000000000000000000000010111111100000000000000000000000: data_out = 6'b110110;
64'b0100000001000000000000000000000010111111100000000000000000000000: data_out = 6'b110111;
64'b0100000010100000000000000000000010111111100000000000000000000000: data_out = 6'b110101;
64'b0100000011100000000000000000000010111111100000000000000000000000: data_out = 6'b110100;
64'b0100000011100000000000000000000011000000010000000000000000000000: data_out = 6'b111100;
64'b0100000010100000000000000000000011000000010000000000000000000000: data_out = 6'b111101;
64'b0100000001000000000000000000000011000000010000000000000000000000: data_out = 6'b111111;
64'b0011111110000000000000000000000011000000010000000000000000000000: data_out = 6'b111110;
64'b1011111110000000000000000000000011000000010000000000000000000000: data_out = 6'b111010;
64'b1100000001000000000000000000000011000000010000000000000000000000: data_out = 6'b111011;
64'b1100000010100000000000000000000011000000010000000000000000000000: data_out = 6'b111001;
64'b1100000011100000000000000000000011000000010000000000000000000000: data_out = 6'b111000;
64'b1100000011100000000000000000000011000000101000000000000000000000: data_out = 6'b101000;
64'b1100000010100000000000000000000011000000101000000000000000000000: data_out = 6'b101001;
64'b1100000001000000000000000000000011000000101000000000000000000000: data_out = 6'b101011;
64'b1011111110000000000000000000000011000000101000000000000000000000: data_out = 6'b101010;
64'b0011111110000000000000000000000011000000101000000000000000000000: data_out = 6'b101110;
64'b0100000001000000000000000000000011000000101000000000000000000000: data_out = 6'b101111;
64'b0100000010100000000000000000000011000000101000000000000000000000: data_out = 6'b101101;
64'b0100000011100000000000000000000011000000101000000000000000000000: data_out = 6'b101100;
64'b0100000011100000000000000000000011000000111000000000000000000000: data_out = 6'b100100;
64'b0100000010100000000000000000000011000000111000000000000000000000: data_out = 6'b100101;
64'b0100000001000000000000000000000011000000111000000000000000000000: data_out = 6'b100111;
64'b0011111110000000000000000000000011000000111000000000000000000000: data_out = 6'b100110;
64'b1011111110000000000000000000000011000000111000000000000000000000: data_out = 6'b100010;
64'b1100000001000000000000000000000011000000111000000000000000000000: data_out = 6'b100011;
64'b1100000010100000000000000000000011000000111000000000000000000000: data_out = 6'b100001;
64'b1100000011100000000000000000000011000000111000000000000000000000: data_out = 6'b100000;
		endcase
	end
endmodule