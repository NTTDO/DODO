module DEQAM_64_imag(
	input [31:0] data_in,
	output reg [5:0] data_out
);
	always@(*)begin
		case(data_in)
			32'b01000000111000000000000000000000: data_out = 6'b000000;
            32'b01000000111000000000000000000000: data_out = 6'b000001;
            32'b01000000111000000000000000000000: data_out = 6'b000011;
            32'b01000000111000000000000000000000: data_out = 6'b000010;
            32'b01000000111000000000000000000000: data_out = 6'b000110;
            32'b01000000111000000000000000000000: data_out = 6'b000111;
            32'b01000000111000000000000000000000: data_out = 6'b000101;
            32'b01000000111000000000000000000000: data_out = 6'b000100;
            32'b01000000101000000000000000000000: data_out = 6'b001100;
            32'b01000000101000000000000000000000: data_out = 6'b001101;
            32'b01000000101000000000000000000000: data_out = 6'b001111;
            32'b01000000101000000000000000000000: data_out = 6'b001110;
            32'b01000000101000000000000000000000: data_out = 6'b001010;
            32'b01000000101000000000000000000000: data_out = 6'b001011;
            32'b01000000101000000000000000000000: data_out = 6'b001001;
            32'b01000000101000000000000000000000: data_out = 6'b001000;
            32'b01000000010000000000000000000000: data_out = 6'b011000;
            32'b01000000010000000000000000000000: data_out = 6'b011001;
            32'b01000000010000000000000000000000: data_out = 6'b011011;
            32'b01000000010000000000000000000000: data_out = 6'b011010;
            32'b01000000010000000000000000000000: data_out = 6'b011110;
            32'b01000000010000000000000000000000: data_out = 6'b011111;
            32'b01000000010000000000000000000000: data_out = 6'b011101;
            32'b01000000010000000000000000000000: data_out = 6'b011100;
            32'b00111111100000000000000000000000: data_out = 6'b010100;
            32'b00111111100000000000000000000000: data_out = 6'b010101;
            32'b00111111100000000000000000000000: data_out = 6'b010111;
            32'b00111111100000000000000000000000: data_out = 6'b010110;
            32'b00111111100000000000000000000000: data_out = 6'b010010;
            32'b00111111100000000000000000000000: data_out = 6'b010011;
            32'b00111111100000000000000000000000: data_out = 6'b010001;
            32'b00111111100000000000000000000000: data_out = 6'b010000;
            32'b10111111100000000000000000000000: data_out = 6'b110000;
            32'b10111111100000000000000000000000: data_out = 6'b110001;
            32'b10111111100000000000000000000000: data_out = 6'b110011;
            32'b10111111100000000000000000000000: data_out = 6'b110010;
            32'b10111111100000000000000000000000: data_out = 6'b110110;
            32'b10111111100000000000000000000000: data_out = 6'b110111;
            32'b10111111100000000000000000000000: data_out = 6'b110101;
            32'b10111111100000000000000000000000: data_out = 6'b110100;
            32'b11000000010000000000000000000000: data_out = 6'b111100;
            32'b11000000010000000000000000000000: data_out = 6'b111101;
            32'b11000000010000000000000000000000: data_out = 6'b111111;
            32'b11000000010000000000000000000000: data_out = 6'b111110;
            32'b11000000010000000000000000000000: data_out = 6'b111010;
            32'b11000000010000000000000000000000: data_out = 6'b111011;
            32'b11000000010000000000000000000000: data_out = 6'b111001;
            32'b11000000010000000000000000000000: data_out = 6'b111000;
            32'b11000000101000000000000000000000: data_out = 6'b101000;
            32'b11000000101000000000000000000000: data_out = 6'b101001;
            32'b11000000101000000000000000000000: data_out = 6'b101011;
            32'b11000000101000000000000000000000: data_out = 6'b101010;
            32'b11000000101000000000000000000000: data_out = 6'b101110;
            32'b11000000101000000000000000000000: data_out = 6'b101111;
            32'b11000000101000000000000000000000: data_out = 6'b101101;
            32'b11000000101000000000000000000000: data_out = 6'b101100;
            32'b11000000111000000000000000000000: data_out = 6'b100100;
            32'b11000000111000000000000000000000: data_out = 6'b100101;
            32'b11000000111000000000000000000000: data_out = 6'b100111;
            32'b11000000111000000000000000000000: data_out = 6'b100110;
            32'b11000000111000000000000000000000: data_out = 6'b100010;
            32'b11000000111000000000000000000000: data_out = 6'b100011;
            32'b11000000111000000000000000000000: data_out = 6'b100001;
            32'b11000000111000000000000000000000: data_out = 6'b100000;
		endcase
	end
endmodule 